-- PRJ_SIM.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PRJ_SIM is
	port (
		AvalonSimpleMaster_0_avm_m0_address     : in    std_logic_vector(7 downto 0)  := (others => '0'); -- AvalonSimpleMaster_0_avm_m0.address
		AvalonSimpleMaster_0_avm_m0_read        : in    std_logic                     := '0';             --                            .read
		AvalonSimpleMaster_0_avm_m0_waitrequest : out   std_logic;                                        --                            .waitrequest
		AvalonSimpleMaster_0_avm_m0_readdata    : out   std_logic_vector(31 downto 0);                    --                            .readdata
		AvalonSimpleMaster_0_avm_m0_write       : in    std_logic                     := '0';             --                            .write
		AvalonSimpleMaster_0_avm_m0_writedata   : in    std_logic_vector(31 downto 0) := (others => '0'); --                            .writedata
		AvalonSimpleMaster_0_reset_reset        : out   std_logic;                                        --  AvalonSimpleMaster_0_reset.reset
		clk_clk                                 : in    std_logic                     := '0';             --                         clk.clk
		pio_0_conduit_end_export                : inout std_logic_vector(7 downto 0)  := (others => '0'); --           pio_0_conduit_end.export
		pio_1_conduit_end_export                : inout std_logic_vector(0 downto 0)  := (others => '0'); --           pio_1_conduit_end.export
		reset_reset_n                           : in    std_logic                     := '0'              --                       reset.reset_n
	);
end entity PRJ_SIM;

architecture rtl of PRJ_SIM is
	component PRJ_SIM_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                          : in  std_logic                     := 'X';             -- clk
			AvalonSimpleMaster_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			AvalonSimpleMaster_0_avm_m0_address                    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			AvalonSimpleMaster_0_avm_m0_waitrequest                : out std_logic;                                        -- waitrequest
			AvalonSimpleMaster_0_avm_m0_read                       : in  std_logic                     := 'X';             -- read
			AvalonSimpleMaster_0_avm_m0_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			AvalonSimpleMaster_0_avm_m0_write                      : in  std_logic                     := 'X';             -- write
			AvalonSimpleMaster_0_avm_m0_writedata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pio_0_avalon_slave_0_address                           : out std_logic_vector(1 downto 0);                     -- address
			pio_0_avalon_slave_0_write                             : out std_logic;                                        -- write
			pio_0_avalon_slave_0_read                              : out std_logic;                                        -- read
			pio_0_avalon_slave_0_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_0_avalon_slave_0_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			pio_0_avalon_slave_0_chipselect                        : out std_logic;                                        -- chipselect
			pio_1_avalon_slave_0_address                           : out std_logic_vector(1 downto 0);                     -- address
			pio_1_avalon_slave_0_write                             : out std_logic;                                        -- write
			pio_1_avalon_slave_0_read                              : out std_logic;                                        -- read
			pio_1_avalon_slave_0_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_1_avalon_slave_0_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			pio_1_avalon_slave_0_chipselect                        : out std_logic                                         -- chipselect
		);
	end component PRJ_SIM_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	component prj_sim_pio_0 is
		generic (
			DATA_WIDTH    : integer := 8;
			PIO_DIRECTION : string  := "OUTPUT"
		);
		port (
			clk          : in    std_logic                     := 'X';             --          clock.clk
			reset_n      : in    std_logic                     := 'X';             --          reset.reset_n
			address      : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- avalon_slave_0.address
			read         : in    std_logic                     := 'X';             --               .read
			readdata     : out   std_logic_vector(31 downto 0);                    --               .readdata
			write        : in    std_logic                     := 'X';             --               .write
			writedata    : in    std_logic_vector(31 downto 0) := (others => 'X'); --               .writedata
			chipselect   : in    std_logic                     := 'X';             --               .chipselect
			pio_external : inout std_logic_vector(7 downto 0)  := (others => 'X')  --    conduit_end.export
		);
	end component prj_sim_pio_0;

	component prj_sim_pio_1 is
		generic (
			DATA_WIDTH    : integer := 8;
			PIO_DIRECTION : string  := "OUTPUT"
		);
		port (
			clk          : in    std_logic                     := 'X';             --          clock.clk
			reset_n      : in    std_logic                     := 'X';             --          reset.reset_n
			address      : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- avalon_slave_0.address
			read         : in    std_logic                     := 'X';             --               .read
			readdata     : out   std_logic_vector(31 downto 0);                    --               .readdata
			write        : in    std_logic                     := 'X';             --               .write
			writedata    : in    std_logic_vector(31 downto 0) := (others => 'X'); --               .writedata
			chipselect   : in    std_logic                     := 'X';             --               .chipselect
			pio_external : inout std_logic_vector(0 downto 0)  := (others => 'X')  --    conduit_end.export
		);
	end component prj_sim_pio_1;

	signal mm_interconnect_0_pio_0_avalon_slave_0_chipselect : std_logic;                     -- mm_interconnect_0:pio_0_avalon_slave_0_chipselect -> pio_0:chipselect
	signal mm_interconnect_0_pio_0_avalon_slave_0_readdata   : std_logic_vector(31 downto 0); -- pio_0:readdata -> mm_interconnect_0:pio_0_avalon_slave_0_readdata
	signal mm_interconnect_0_pio_0_avalon_slave_0_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_0_avalon_slave_0_address -> pio_0:address
	signal mm_interconnect_0_pio_0_avalon_slave_0_read       : std_logic;                     -- mm_interconnect_0:pio_0_avalon_slave_0_read -> pio_0:read
	signal mm_interconnect_0_pio_0_avalon_slave_0_write      : std_logic;                     -- mm_interconnect_0:pio_0_avalon_slave_0_write -> pio_0:write
	signal mm_interconnect_0_pio_0_avalon_slave_0_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_0_avalon_slave_0_writedata -> pio_0:writedata
	signal mm_interconnect_0_pio_1_avalon_slave_0_chipselect : std_logic;                     -- mm_interconnect_0:pio_1_avalon_slave_0_chipselect -> pio_1:chipselect
	signal mm_interconnect_0_pio_1_avalon_slave_0_readdata   : std_logic_vector(31 downto 0); -- pio_1:readdata -> mm_interconnect_0:pio_1_avalon_slave_0_readdata
	signal mm_interconnect_0_pio_1_avalon_slave_0_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_1_avalon_slave_0_address -> pio_1:address
	signal mm_interconnect_0_pio_1_avalon_slave_0_read       : std_logic;                     -- mm_interconnect_0:pio_1_avalon_slave_0_read -> pio_1:read
	signal mm_interconnect_0_pio_1_avalon_slave_0_write      : std_logic;                     -- mm_interconnect_0:pio_1_avalon_slave_0_write -> pio_1:write
	signal mm_interconnect_0_pio_1_avalon_slave_0_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_1_avalon_slave_0_writedata -> pio_1:writedata
	signal rst_controller_reset_out_reset                    : std_logic;                     -- rst_controller:reset_out -> [AvalonSimpleMaster_0_reset_reset, AvalonSimpleMaster_0_reset_reset:in, mm_interconnect_0:AvalonSimpleMaster_0_reset_reset_bridge_in_reset_reset]
	signal reset_reset_n_ports_inv                           : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal avalonsimplemaster_0_reset_reset_ports_inv        : std_logic;                     -- AvalonSimpleMaster_0_reset_reset:inv -> [pio_0:reset_n, pio_1:reset_n]

begin

	pio_0 : component prj_sim_pio_0
		generic map (
			DATA_WIDTH    => 8,
			PIO_DIRECTION => "OUTPUT"
		)
		port map (
			clk          => clk_clk,                                           --          clock.clk
			reset_n      => avalonsimplemaster_0_reset_reset_ports_inv,        --          reset.reset_n
			address      => mm_interconnect_0_pio_0_avalon_slave_0_address,    -- avalon_slave_0.address
			read         => mm_interconnect_0_pio_0_avalon_slave_0_read,       --               .read
			readdata     => mm_interconnect_0_pio_0_avalon_slave_0_readdata,   --               .readdata
			write        => mm_interconnect_0_pio_0_avalon_slave_0_write,      --               .write
			writedata    => mm_interconnect_0_pio_0_avalon_slave_0_writedata,  --               .writedata
			chipselect   => mm_interconnect_0_pio_0_avalon_slave_0_chipselect, --               .chipselect
			pio_external => pio_0_conduit_end_export                           --    conduit_end.export
		);

	pio_1 : component prj_sim_pio_1
		generic map (
			DATA_WIDTH    => 1,
			PIO_DIRECTION => "INPUT"
		)
		port map (
			clk          => clk_clk,                                           --          clock.clk
			reset_n      => avalonsimplemaster_0_reset_reset_ports_inv,        --          reset.reset_n
			address      => mm_interconnect_0_pio_1_avalon_slave_0_address,    -- avalon_slave_0.address
			read         => mm_interconnect_0_pio_1_avalon_slave_0_read,       --               .read
			readdata     => mm_interconnect_0_pio_1_avalon_slave_0_readdata,   --               .readdata
			write        => mm_interconnect_0_pio_1_avalon_slave_0_write,      --               .write
			writedata    => mm_interconnect_0_pio_1_avalon_slave_0_writedata,  --               .writedata
			chipselect   => mm_interconnect_0_pio_1_avalon_slave_0_chipselect, --               .chipselect
			pio_external => pio_1_conduit_end_export                           --    conduit_end.export
		);

	mm_interconnect_0 : component PRJ_SIM_mm_interconnect_0
		port map (
			clk_0_clk_clk                                          => clk_clk,                                           --                                        clk_0_clk.clk
			AvalonSimpleMaster_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                    -- AvalonSimpleMaster_0_reset_reset_bridge_in_reset.reset
			AvalonSimpleMaster_0_avm_m0_address                    => AvalonSimpleMaster_0_avm_m0_address,               --                      AvalonSimpleMaster_0_avm_m0.address
			AvalonSimpleMaster_0_avm_m0_waitrequest                => AvalonSimpleMaster_0_avm_m0_waitrequest,           --                                                 .waitrequest
			AvalonSimpleMaster_0_avm_m0_read                       => AvalonSimpleMaster_0_avm_m0_read,                  --                                                 .read
			AvalonSimpleMaster_0_avm_m0_readdata                   => AvalonSimpleMaster_0_avm_m0_readdata,              --                                                 .readdata
			AvalonSimpleMaster_0_avm_m0_write                      => AvalonSimpleMaster_0_avm_m0_write,                 --                                                 .write
			AvalonSimpleMaster_0_avm_m0_writedata                  => AvalonSimpleMaster_0_avm_m0_writedata,             --                                                 .writedata
			pio_0_avalon_slave_0_address                           => mm_interconnect_0_pio_0_avalon_slave_0_address,    --                             pio_0_avalon_slave_0.address
			pio_0_avalon_slave_0_write                             => mm_interconnect_0_pio_0_avalon_slave_0_write,      --                                                 .write
			pio_0_avalon_slave_0_read                              => mm_interconnect_0_pio_0_avalon_slave_0_read,       --                                                 .read
			pio_0_avalon_slave_0_readdata                          => mm_interconnect_0_pio_0_avalon_slave_0_readdata,   --                                                 .readdata
			pio_0_avalon_slave_0_writedata                         => mm_interconnect_0_pio_0_avalon_slave_0_writedata,  --                                                 .writedata
			pio_0_avalon_slave_0_chipselect                        => mm_interconnect_0_pio_0_avalon_slave_0_chipselect, --                                                 .chipselect
			pio_1_avalon_slave_0_address                           => mm_interconnect_0_pio_1_avalon_slave_0_address,    --                             pio_1_avalon_slave_0.address
			pio_1_avalon_slave_0_write                             => mm_interconnect_0_pio_1_avalon_slave_0_write,      --                                                 .write
			pio_1_avalon_slave_0_read                              => mm_interconnect_0_pio_1_avalon_slave_0_read,       --                                                 .read
			pio_1_avalon_slave_0_readdata                          => mm_interconnect_0_pio_1_avalon_slave_0_readdata,   --                                                 .readdata
			pio_1_avalon_slave_0_writedata                         => mm_interconnect_0_pio_1_avalon_slave_0_writedata,  --                                                 .writedata
			pio_1_avalon_slave_0_chipselect                        => mm_interconnect_0_pio_1_avalon_slave_0_chipselect  --                                                 .chipselect
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	avalonsimplemaster_0_reset_reset_ports_inv <= not rst_controller_reset_out_reset;

	AvalonSimpleMaster_0_reset_reset <= rst_controller_reset_out_reset;

end architecture rtl; -- of PRJ_SIM
