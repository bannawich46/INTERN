
module Assignment4 (
	clk_clk,
	reset_reset_n,
	pio_0_conduit_end_export);	

	input		clk_clk;
	input		reset_reset_n;
	inout	[8:0]	pio_0_conduit_end_export;
endmodule
