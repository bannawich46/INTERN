
module Assignment5 (
	clk_clk,
	reset_reset_n,
	pwm_0_conduit_end_writedata);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	pwm_0_conduit_end_writedata;
endmodule
