-- PRJ_SIM.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PRJ_SIM is
	port (
		Avalon_Simple_Master_0_avm_m0_address     : in  std_logic_vector(8 downto 0)  := (others => '0'); -- Avalon_Simple_Master_0_avm_m0.address
		Avalon_Simple_Master_0_avm_m0_read        : in  std_logic                     := '0';             --                              .read
		Avalon_Simple_Master_0_avm_m0_waitrequest : out std_logic;                                        --                              .waitrequest
		Avalon_Simple_Master_0_avm_m0_readdata    : out std_logic_vector(31 downto 0);                    --                              .readdata
		Avalon_Simple_Master_0_avm_m0_write       : in  std_logic                     := '0';             --                              .write
		Avalon_Simple_Master_0_avm_m0_writedata   : in  std_logic_vector(31 downto 0) := (others => '0'); --                              .writedata
		Avalon_Simple_Master_0_reset_reset        : out std_logic;                                        --  Avalon_Simple_Master_0_reset.reset
		clk_clk                                   : in  std_logic                     := '0';             --                           clk.clk
		ocram_master_0_conduit_end_export         : out std_logic_vector(7 downto 0);                     --    ocram_master_0_conduit_end.export
		reset_reset_n                             : in  std_logic                     := '0'              --                         reset.reset_n
	);
end entity PRJ_SIM;

architecture rtl of PRJ_SIM is
	component OCRAM_MASTER is
		port (
			CLK                : in  std_logic                     := 'X';             -- clk
			iADDRESS           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			iREAD              : in  std_logic                     := 'X';             -- read
			iREADDATA          : out std_logic_vector(31 downto 0);                    -- readdata
			iCHIPSELECT        : in  std_logic                     := 'X';             -- chipselect
			iWAITREQUEST       : out std_logic;                                        -- waitrequest
			iADDRESS_OCRAM     : out std_logic_vector(9 downto 0);                     -- address
			iREADDATA_OCRAM    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			iREAD_OCRAM        : out std_logic;                                        -- read
			iWAITREQUEST_OCRAM : in  std_logic                     := 'X';             -- waitrequest
			RST                : in  std_logic                     := 'X';             -- reset
			EXTERNAL           : out std_logic_vector(7 downto 0)                      -- export
		);
	end component OCRAM_MASTER;

	component PRJ_SIM_onchip_memory2_0 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component PRJ_SIM_onchip_memory2_0;

	component PRJ_SIM_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                         : in  std_logic                     := 'X';             -- clk
			ocram_master_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			ocram_master_0_avalon_master_address                  : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			ocram_master_0_avalon_master_waitrequest              : out std_logic;                                        -- waitrequest
			ocram_master_0_avalon_master_read                     : in  std_logic                     := 'X';             -- read
			ocram_master_0_avalon_master_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			onchip_memory2_0_s2_address                           : out std_logic_vector(5 downto 0);                     -- address
			onchip_memory2_0_s2_write                             : out std_logic;                                        -- write
			onchip_memory2_0_s2_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s2_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s2_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s2_chipselect                        : out std_logic;                                        -- chipselect
			onchip_memory2_0_s2_clken                             : out std_logic                                         -- clken
		);
	end component PRJ_SIM_mm_interconnect_0;

	component PRJ_SIM_mm_interconnect_1 is
		port (
			clk_0_clk_clk                                            : in  std_logic                     := 'X';             -- clk
			Avalon_Simple_Master_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Avalon_Simple_Master_0_avm_m0_address                    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			Avalon_Simple_Master_0_avm_m0_waitrequest                : out std_logic;                                        -- waitrequest
			Avalon_Simple_Master_0_avm_m0_read                       : in  std_logic                     := 'X';             -- read
			Avalon_Simple_Master_0_avm_m0_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			Avalon_Simple_Master_0_avm_m0_write                      : in  std_logic                     := 'X';             -- write
			Avalon_Simple_Master_0_avm_m0_writedata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			ocram_master_0_avalon_slave_0_address                    : out std_logic_vector(1 downto 0);                     -- address
			ocram_master_0_avalon_slave_0_read                       : out std_logic;                                        -- read
			ocram_master_0_avalon_slave_0_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ocram_master_0_avalon_slave_0_waitrequest                : in  std_logic                     := 'X';             -- waitrequest
			ocram_master_0_avalon_slave_0_chipselect                 : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_address                              : out std_logic_vector(5 downto 0);                     -- address
			onchip_memory2_0_s1_write                                : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                           : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                           : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                                : out std_logic                                         -- clken
		);
	end component PRJ_SIM_mm_interconnect_1;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal ocram_master_0_avalon_master_readdata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:ocram_master_0_avalon_master_readdata -> ocram_master_0:iREADDATA_OCRAM
	signal ocram_master_0_avalon_master_waitrequest                    : std_logic;                     -- mm_interconnect_0:ocram_master_0_avalon_master_waitrequest -> ocram_master_0:iWAITREQUEST_OCRAM
	signal ocram_master_0_avalon_master_address                        : std_logic_vector(9 downto 0);  -- ocram_master_0:iADDRESS_OCRAM -> mm_interconnect_0:ocram_master_0_avalon_master_address
	signal ocram_master_0_avalon_master_read                           : std_logic;                     -- ocram_master_0:iREAD_OCRAM -> mm_interconnect_0:ocram_master_0_avalon_master_read
	signal mm_interconnect_0_onchip_memory2_0_s2_chipselect            : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	signal mm_interconnect_0_onchip_memory2_0_s2_readdata              : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata2 -> mm_interconnect_0:onchip_memory2_0_s2_readdata
	signal mm_interconnect_0_onchip_memory2_0_s2_address               : std_logic_vector(5 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	signal mm_interconnect_0_onchip_memory2_0_s2_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s2_byteenable -> onchip_memory2_0:byteenable2
	signal mm_interconnect_0_onchip_memory2_0_s2_write                 : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	signal mm_interconnect_0_onchip_memory2_0_s2_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	signal mm_interconnect_0_onchip_memory2_0_s2_clken                 : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	signal mm_interconnect_1_ocram_master_0_avalon_slave_0_chipselect  : std_logic;                     -- mm_interconnect_1:ocram_master_0_avalon_slave_0_chipselect -> ocram_master_0:iCHIPSELECT
	signal mm_interconnect_1_ocram_master_0_avalon_slave_0_readdata    : std_logic_vector(31 downto 0); -- ocram_master_0:iREADDATA -> mm_interconnect_1:ocram_master_0_avalon_slave_0_readdata
	signal mm_interconnect_1_ocram_master_0_avalon_slave_0_waitrequest : std_logic;                     -- ocram_master_0:iWAITREQUEST -> mm_interconnect_1:ocram_master_0_avalon_slave_0_waitrequest
	signal mm_interconnect_1_ocram_master_0_avalon_slave_0_address     : std_logic_vector(1 downto 0);  -- mm_interconnect_1:ocram_master_0_avalon_slave_0_address -> ocram_master_0:iADDRESS
	signal mm_interconnect_1_ocram_master_0_avalon_slave_0_read        : std_logic;                     -- mm_interconnect_1:ocram_master_0_avalon_slave_0_read -> ocram_master_0:iREAD
	signal mm_interconnect_1_onchip_memory2_0_s1_chipselect            : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_1_onchip_memory2_0_s1_readdata              : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_1:onchip_memory2_0_s1_readdata
	signal mm_interconnect_1_onchip_memory2_0_s1_address               : std_logic_vector(5 downto 0);  -- mm_interconnect_1:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_1_onchip_memory2_0_s1_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_1:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_1_onchip_memory2_0_s1_write                 : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_1_onchip_memory2_0_s1_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_1:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_1_onchip_memory2_0_s1_clken                 : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal rst_controller_reset_out_reset                              : std_logic;                     -- rst_controller:reset_out -> [Avalon_Simple_Master_0_reset_reset, mm_interconnect_0:ocram_master_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:Avalon_Simple_Master_0_reset_reset_bridge_in_reset_reset, ocram_master_0:RST, onchip_memory2_0:reset, onchip_memory2_0:reset2, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                          : std_logic;                     -- rst_controller:reset_req -> [onchip_memory2_0:reset_req, onchip_memory2_0:reset_req2, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                     : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0

begin

	ocram_master_0 : component OCRAM_MASTER
		port map (
			CLK                => clk_clk,                                                     --          clock.clk
			iADDRESS           => mm_interconnect_1_ocram_master_0_avalon_slave_0_address,     -- avalon_slave_0.address
			iREAD              => mm_interconnect_1_ocram_master_0_avalon_slave_0_read,        --               .read
			iREADDATA          => mm_interconnect_1_ocram_master_0_avalon_slave_0_readdata,    --               .readdata
			iCHIPSELECT        => mm_interconnect_1_ocram_master_0_avalon_slave_0_chipselect,  --               .chipselect
			iWAITREQUEST       => mm_interconnect_1_ocram_master_0_avalon_slave_0_waitrequest, --               .waitrequest
			iADDRESS_OCRAM     => ocram_master_0_avalon_master_address,                        --  avalon_master.address
			iREADDATA_OCRAM    => ocram_master_0_avalon_master_readdata,                       --               .readdata
			iREAD_OCRAM        => ocram_master_0_avalon_master_read,                           --               .read
			iWAITREQUEST_OCRAM => ocram_master_0_avalon_master_waitrequest,                    --               .waitrequest
			RST                => rst_controller_reset_out_reset,                              --     reset_sink.reset
			EXTERNAL           => ocram_master_0_conduit_end_export                            --    conduit_end.export
		);

	onchip_memory2_0 : component PRJ_SIM_onchip_memory2_0
		port map (
			clk         => clk_clk,                                          --   clk1.clk
			address     => mm_interconnect_1_onchip_memory2_0_s1_address,    --     s1.address
			clken       => mm_interconnect_1_onchip_memory2_0_s1_clken,      --       .clken
			chipselect  => mm_interconnect_1_onchip_memory2_0_s1_chipselect, --       .chipselect
			write       => mm_interconnect_1_onchip_memory2_0_s1_write,      --       .write
			readdata    => mm_interconnect_1_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_1_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_1_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,               --       .reset_req
			address2    => mm_interconnect_0_onchip_memory2_0_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_onchip_memory2_0_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_onchip_memory2_0_s2_clken,      --       .clken
			write2      => mm_interconnect_0_onchip_memory2_0_s2_write,      --       .write
			readdata2   => mm_interconnect_0_onchip_memory2_0_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_onchip_memory2_0_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_onchip_memory2_0_s2_byteenable, --       .byteenable
			clk2        => clk_clk,                                          --   clk2.clk
			reset2      => rst_controller_reset_out_reset,                   -- reset2.reset
			reset_req2  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze      => '0'                                               -- (terminated)
		);

	mm_interconnect_0 : component PRJ_SIM_mm_interconnect_0
		port map (
			clk_0_clk_clk                                         => clk_clk,                                          --                                       clk_0_clk.clk
			ocram_master_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                   -- ocram_master_0_reset_sink_reset_bridge_in_reset.reset
			ocram_master_0_avalon_master_address                  => ocram_master_0_avalon_master_address,             --                    ocram_master_0_avalon_master.address
			ocram_master_0_avalon_master_waitrequest              => ocram_master_0_avalon_master_waitrequest,         --                                                .waitrequest
			ocram_master_0_avalon_master_read                     => ocram_master_0_avalon_master_read,                --                                                .read
			ocram_master_0_avalon_master_readdata                 => ocram_master_0_avalon_master_readdata,            --                                                .readdata
			onchip_memory2_0_s2_address                           => mm_interconnect_0_onchip_memory2_0_s2_address,    --                             onchip_memory2_0_s2.address
			onchip_memory2_0_s2_write                             => mm_interconnect_0_onchip_memory2_0_s2_write,      --                                                .write
			onchip_memory2_0_s2_readdata                          => mm_interconnect_0_onchip_memory2_0_s2_readdata,   --                                                .readdata
			onchip_memory2_0_s2_writedata                         => mm_interconnect_0_onchip_memory2_0_s2_writedata,  --                                                .writedata
			onchip_memory2_0_s2_byteenable                        => mm_interconnect_0_onchip_memory2_0_s2_byteenable, --                                                .byteenable
			onchip_memory2_0_s2_chipselect                        => mm_interconnect_0_onchip_memory2_0_s2_chipselect, --                                                .chipselect
			onchip_memory2_0_s2_clken                             => mm_interconnect_0_onchip_memory2_0_s2_clken       --                                                .clken
		);

	mm_interconnect_1 : component PRJ_SIM_mm_interconnect_1
		port map (
			clk_0_clk_clk                                            => clk_clk,                                                     --                                          clk_0_clk.clk
			Avalon_Simple_Master_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                              -- Avalon_Simple_Master_0_reset_reset_bridge_in_reset.reset
			Avalon_Simple_Master_0_avm_m0_address                    => Avalon_Simple_Master_0_avm_m0_address,                       --                      Avalon_Simple_Master_0_avm_m0.address
			Avalon_Simple_Master_0_avm_m0_waitrequest                => Avalon_Simple_Master_0_avm_m0_waitrequest,                   --                                                   .waitrequest
			Avalon_Simple_Master_0_avm_m0_read                       => Avalon_Simple_Master_0_avm_m0_read,                          --                                                   .read
			Avalon_Simple_Master_0_avm_m0_readdata                   => Avalon_Simple_Master_0_avm_m0_readdata,                      --                                                   .readdata
			Avalon_Simple_Master_0_avm_m0_write                      => Avalon_Simple_Master_0_avm_m0_write,                         --                                                   .write
			Avalon_Simple_Master_0_avm_m0_writedata                  => Avalon_Simple_Master_0_avm_m0_writedata,                     --                                                   .writedata
			ocram_master_0_avalon_slave_0_address                    => mm_interconnect_1_ocram_master_0_avalon_slave_0_address,     --                      ocram_master_0_avalon_slave_0.address
			ocram_master_0_avalon_slave_0_read                       => mm_interconnect_1_ocram_master_0_avalon_slave_0_read,        --                                                   .read
			ocram_master_0_avalon_slave_0_readdata                   => mm_interconnect_1_ocram_master_0_avalon_slave_0_readdata,    --                                                   .readdata
			ocram_master_0_avalon_slave_0_waitrequest                => mm_interconnect_1_ocram_master_0_avalon_slave_0_waitrequest, --                                                   .waitrequest
			ocram_master_0_avalon_slave_0_chipselect                 => mm_interconnect_1_ocram_master_0_avalon_slave_0_chipselect,  --                                                   .chipselect
			onchip_memory2_0_s1_address                              => mm_interconnect_1_onchip_memory2_0_s1_address,               --                                onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                                => mm_interconnect_1_onchip_memory2_0_s1_write,                 --                                                   .write
			onchip_memory2_0_s1_readdata                             => mm_interconnect_1_onchip_memory2_0_s1_readdata,              --                                                   .readdata
			onchip_memory2_0_s1_writedata                            => mm_interconnect_1_onchip_memory2_0_s1_writedata,             --                                                   .writedata
			onchip_memory2_0_s1_byteenable                           => mm_interconnect_1_onchip_memory2_0_s1_byteenable,            --                                                   .byteenable
			onchip_memory2_0_s1_chipselect                           => mm_interconnect_1_onchip_memory2_0_s1_chipselect,            --                                                   .chipselect
			onchip_memory2_0_s1_clken                                => mm_interconnect_1_onchip_memory2_0_s1_clken                  --                                                   .clken
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	Avalon_Simple_Master_0_reset_reset <= rst_controller_reset_out_reset;

end architecture rtl; -- of PRJ_SIM
